`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:42:02 09/20/2017 
// Design Name: 
// Module Name:    vga_r 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vga_r(
    output reg red,
    output reg green,
    output reg blue,
    input [9:0] pos_h,
    input [9:0] pos_v,
    input blank,
    input clk,
    input SW0,
    input SW1,
    input SW2
    );


endmodule
