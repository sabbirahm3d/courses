`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:53:16 10/09/2017 
// Design Name: 
// Module Name:    igniter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module igniter(
		output position,
		input [3:0] delta,
		input enable_jump,
		input sys_clk,
		input clr_n
	);




endmodule
